`define STATUS          12
`define CAUSE           13
`define EPC             14
`define SYSCALL   5'b01000
`define BREAK     5'b01001
`define TEQ       5'b01101

`define ADD_op          6'b000000
`define SUB_op          6'b000000
`define ADDU_op         6'b000000
`define SUBU_op         6'b000000
`define AND_op          6'b000000
`define JR_op           6'b000000
`define XOR_op          6'b000000
`define NOR_op          6'b000000
`define OR_op           6'b000000
`define SLT_op          6'b000000
`define SRLV_op         6'b000000
`define SRAV_op         6'b000000
`define SLL_op          6'b000000
`define SLLV_op         6'b000000
`define SLTU_op         6'b000000
`define SRA_op          6'b000000
`define SRL_op          6'b000000
`define ADDI_op         6'b001000
`define ADDIU_op        6'b001001
`define ANDI_op         6'b001100
`define ORI_op          6'b001101
`define SLTIU_op        6'b001011
`define LUI_op          6'b001111
`define XORI_op         6'b001110
`define SLTI_op         6'b001010
`define SW_op           6'b101011
`define LW_op           6'b100011
`define BEQ_op          6'b000100
`define BNE_op          6'b000101
`define CLZ_op          6'b011100
`define DIVU_op         6'b000000
`define ERET_op         6'b010000
`define LHU_op          6'b100101
`define SB_op           6'b101000
`define SH_op           6'b101001
`define LH_op           6'b100001
`define MFHI_op         6'b000000
`define MFLO_op         6'b000000
`define MTHI_op         6'b000000
`define MTLO_op         6'b000000
`define MUL_op          6'b011100
`define MULTU_op        6'b000000
`define SYSCALL_op      6'b000000
`define TEQ_op          6'b000000
`define BGEZ_op         6'b000001
`define BREAK_op        6'b000000
`define DIV_op          6'b000000
`define J_op            6'b000010
`define JAL_op          6'b000011
`define JALR_op         6'b000000
`define LB_op           6'b100000
`define LBU_op          6'b100100


`define ADD_func        6'b100000
`define SUB_func        6'b100010
`define ADDU_func       6'b100001
`define SUBU_func       6'b100011
`define AND_func        6'b100100
`define XOR_func        6'b100110
`define NOR_func        6'b100111
`define OR_func         6'b100101
`define SLL_func        6'b000000
`define SLLV_func       6'b000100
`define SLTU_func       6'b101011
`define SRA_func        6'b000011
`define SRL_func        6'b000010
`define SLT_func        6'b101010
`define SRLV_func       6'b000110
`define SRAV_func       6'b000111
`define JR_func         6'b001000
`define CLZ_func        6'b100000
`define DIVU_func       6'b011011
`define ERET_func       6'b011000
`define JALR_func       6'b001001
`define MFHI_func       6'b010000
`define MFLO_func       6'b010010
`define MTHI_func       6'b010001
`define MTLO_func       6'b010011
`define MUL_func        6'b000010
`define MULTU_func      6'b011001
`define SYSCALL_func    6'b001100
`define TEQ_func        6'b110100
`define BREAK_func      6'b001101
`define DIV_func        6'b011010
